-------------------------------------------------------------------------------
--
-- Module Name: prog_mem
-- Create Date: 11/30/2014
-- Description: 
--
-------------------------------------------------------------------------------